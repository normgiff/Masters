** Profile: "SCHEMATIC1-run1"  [ C:\Users\dkhoury\Desktop\SourceTree-Masters\explorations\power\AdjustableVoltageRegulator-PSpiceFiles\SCHEMATIC1\run1.sim ] 

** Creating circuit file "run1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/dkhoury/OneDrive/Documents/pspice_libraries/opamp.lib" 
.LIB "C:/Users/dkhoury/OneDrive/Documents/pspice_libraries/diode.lib" 
* From [PSPICE NETLIST] section of C:\Users\dkhoury\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
