`timescale 1ns / 1ps

// Top Verilog module.
module TOP_MODULE(CLK, RST, OUTPUT_SIG);
	input CLK;
	input RST; 
	
	output [127:0] OUTPUT_SIG;
	

endmodule
