`timescale 1ns / 1ps

module CENTRAL_FSM(
    );


endmodule
