`timescale 1ns / 1ps

/* 
 * Author: Daniel Khoury
 *
 * Generates random values from a seed using a LFSR (linear feedback shift register) circuit.
 */
module RANDOM_GEN(CLK, RST, LOAD_SEED, GET_NEXT, SEED, VAL);
	input CLK;
	input RST;
	input LOAD_SEED;
	input GET_NEXT;
	input [7:0] SEED;
	
	output [7:0] VAL;
	
	LFSR LFSR_ARR0 (.CLK(CLK), .RST(RST), .SEED(SEED[3:0]), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[0]));
	LFSR LFSR_ARR1 (.CLK(CLK), .RST(RST), .SEED(SEED[4:1]), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[1]));
	LFSR LFSR_ARR2 (.CLK(CLK), .RST(RST), .SEED(SEED[5:2]), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[2]));
	LFSR LFSR_ARR3 (.CLK(CLK), .RST(RST), .SEED(SEED[6:3]), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[3]));
	LFSR LFSR_ARR4 (.CLK(CLK), .RST(RST), .SEED(SEED[7:4]), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[4]));
	LFSR LFSR_ARR5 (.CLK(CLK), .RST(RST), .SEED({SEED[2], SEED[0], SEED[5], SEED[1]}), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[5]));
	LFSR LFSR_ARR6 (.CLK(CLK), .RST(RST), .SEED({SEED[5], SEED[3], SEED[7], SEED[6]}), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[6]));
	LFSR LFSR_ARR7 (.CLK(CLK), .RST(RST), .SEED({SEED[0], SEED[3], SEED[4], SEED[7]}), .LOAD(LOAD_SEED), .GET_NEXT(GET_NEXT), .OUT(VAL[7]));
	
endmodule
